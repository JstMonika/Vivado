`timescale 1ns/1ps

module Mux_1bit (a, b, sel, f);
input a, b;
input sel;
output f;

endmodule
