`timescale 1ns/1ps

module FullAdder (a, b, cin, cout, sum);
input a, b;
input cin;
output sum;
output cout;

endmodule
